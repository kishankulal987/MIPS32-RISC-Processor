module adder(input [31:0]A,output [31:0]out);
assign out=A+1'b1;
endmodule